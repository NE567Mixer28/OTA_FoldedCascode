** sch_path: /home/ttuser/OTA_FoldedCascode/xschem/Polarizzazione_Pmos.sch
**.subckt Polarizzazione_Pmos
V1 GND G 1.1
V2 GND D 1.8
XM1 D G GND GND sky130_fd_pr__pfet_01v8 L=2 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code



* ngspice commands

.options savecurrents
*.dc v2 0 1.8 0.01
.control
save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
op
remzerovec
write Polarizzazione_Pmos.raw

.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
